
MACRO "serpentine_50px_0
  CLASS CORE ;
  ORIGIN  0 0 ;
  FOREIGN "serpentine_50px_0 0 0 ;
  SIZE 300 BY 300 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN fl_in1
    DIRECTION 1 ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.5 29.5 30.5 30.5 ;
    END
  END fl_in1
  PIN fl_out
    DIRECTION 1 ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 32.5 32.5 34.5 34.5 ;
    END
  END fl_out
  PIN fl_in2
    DIRECTION 1 ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 36.5 36.5 38.5 38.5 ;
    END
  END fl_in2
  OBS
    LAYER met1 ;
      RECT 0 300.5 0 300.6 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END "serpentine_50px_0