
MACRO %Name%
  CLASS CORE ;
  ORIGIN  %Org_1X% %Org_1Y% ;
  FOREIGN %Name% 0 0 ;
  SIZE %Bounds.x% BY %Bounds.y% ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN %Pin_#[%
    DIRECTION %Pin_#.Dir% ;
    USE SIGNAL ;
    PORT
      LAYER %Pin_#.Layer% ;
        RECT %Pin_#.X1% %Pin_#.Y1% %Pin_#.X2% %Pin_#.Y2% ;
    END
  END %Pin_#]%
  OBS
    LAYER %OBS.Layer% ;
      RECT %OBS.X1% %OBS.Y1% %OBS.X2% %OBS.Y2% ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END %Name%